library verilog;
use verilog.vl_types.all;
entity ALU_Test_vlg_vec_tst is
end ALU_Test_vlg_vec_tst;
