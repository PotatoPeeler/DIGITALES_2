library verilog;
use verilog.vl_types.all;
entity Memory_Test_vlg_vec_tst is
end Memory_Test_vlg_vec_tst;
