library verilog;
use verilog.vl_types.all;
entity Half_adder_vlg_vec_tst is
end Half_adder_vlg_vec_tst;
