library verilog;
use verilog.vl_types.all;
entity MemoriaROM_vlg_vec_tst is
end MemoriaROM_vlg_vec_tst;
