library verilog;
use verilog.vl_types.all;
entity Outputs_Ports1_vlg_vec_tst is
end Outputs_Ports1_vlg_vec_tst;
