library verilog;
use verilog.vl_types.all;
entity DECO_HEX_vlg_vec_tst is
end DECO_HEX_vlg_vec_tst;
