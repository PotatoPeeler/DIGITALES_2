library verilog;
use verilog.vl_types.all;
entity Deco_7Seg_vlg_vec_tst is
end Deco_7Seg_vlg_vec_tst;
