library verilog;
use verilog.vl_types.all;
entity RAM_16x8_sync_vlg_vec_tst is
end RAM_16x8_sync_vlg_vec_tst;
